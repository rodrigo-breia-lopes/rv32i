//module top (
//    input wire clk,
//    input wire rst,
//    input wire read,
//    input wire data,
//    output 
//
//);
//    
//endmodule
